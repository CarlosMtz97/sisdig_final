----------------------------------------------------------------------------------
-- Company:        
-- Engineer:       
-- 
-- Create Date:    
-- Design Name: 
-- Module Name:    VGA_DISPLAY - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description:    
--  
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
-- Commonly used libraries
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity VGA_DISPLAY is
  Generic
  ( n         : integer := 14;                    -- Number of Address bus lines, for an image of 128x128 pixels
	 m         : integer := 8);                    -- Number of Data bus lines
  port (
	 Xin       : in  STD_LOGIC_VECTOR(9 downto 0); -- Column screen coordinate
	 Yin       : in  STD_LOGIC_VECTOR(9 downto 0); -- Row screen coordinate
	 En        : in  STD_LOGIC;                    -- When '1', pixels can be drawn 
	 Enable60  : in  STD_LOGIC;                    -- Enable for cookie
	 rightB    : in  STD_LOGIC;                    -- Right button
	 leftB     : in  STD_LOGIC;                    -- Left button
	 rst       : in  STD_LOGIC;                    -- Reset
	 clk       : in  STD_LOGIC;                    -- Clock from FPGA
	 R   		  : out STD_LOGIC_VECTOR(2 downto 0); -- 3-bit Red channel
	 G   		  : out STD_LOGIC_VECTOR(2 downto 0); -- 3-bit Green channel
	 B   		  : out STD_LOGIC_VECTOR(1 downto 0));-- 2-bit Blue channel
end VGA_DISPLAY;


architecture Behavioral of VGA_DISPLAY is
  -- Embedded signal to group the colors into 1-byte
  -- The colors will be as follows:
  --  R2 R1 R0 G2 G1 G0 B1 B0
  signal Color        : STD_LOGIC_VECTOR(7 downto 0); 
  signal Color_Cookie : STD_LOGIC_VECTOR(7 downto 0); 
  
  --Addresses for the different images that will be displayed
  signal AddressCookie       : STD_LOGIC_VECTOR(n-1 downto 0);  --Super Cookie
  signal AddressCookieL      : STD_LOGIC_VECTOR(n-1 downto 0);  --Super Cookie Left
  signal AddressCookieR      : STD_LOGIC_VECTOR(n-1 downto 0);  --Super Cookie Right
  signal Data              : STD_LOGIC_VECTOR(m-1 downto 0);
  
  --Types of roms that will be used
  type characterImage is array (0 to (128**2) - 1) of STD_LOGIC_VECTOR (7 downto 0);
 
  constant cookieF : characterImage := (
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FB",x"B2",x"8D",
x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"89",x"B1",x"DB",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"D6",x"8D",x"64",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"68",x"B2",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"DA",x"68",x"44",x"44",x"44",x"64",x"68",
x"88",x"8C",x"AC",x"AC",x"AD",x"AC",x"AC",x"AC",x"88",x"68",x"64",x"44",x"44",x"44",x"68",x"B2",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"8D",x"64",x"44",x"64",x"68",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"88",x"64",x"44",x"44",
x"68",x"DA",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",x"68",x"44",x"64",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"64",
x"44",x"64",x"B1",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"64",x"44",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"88",x"64",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"B2",x"64",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"64",x"44",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"B2",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"64",x"44",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"B6",x"64",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"89",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"DA",x"64",x"64",x"B1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",
x"F6",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"68",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",
x"FB",x"D1",x"D1",x"D1",x"D1",x"B1",x"64",x"44",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",
x"8D",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",
x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"64",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",
x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D5",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",
x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"F5",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FA",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",
x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"F5",x"FF",x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"D5",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"68",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",
x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"FF",x"FF",x"FA",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"64",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",
x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"68",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"68",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",
x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"D5",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"DB",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"AC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"8D",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"64",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"68",x"FF",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"68",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FA",x"D5",x"FF",
x"FF",x"FB",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F5",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"DA",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FA",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"FF",
x"FF",x"FA",x"D5",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"F6",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B1",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"91",x"44",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D5",x"FA",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"FA",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"44",x"89",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"64",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",
x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"68",x"D1",x"D1",x"D5",
x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"FA",x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",
x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"DB",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"44",x"88",x"D1",x"FB",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FA",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",
x"FF",x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"D6",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"8C",x"D1",x"FB",x"FF",
x"FB",x"FA",x"D5",x"D1",x"D1",x"D1",x"D5",x"F6",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"DF",
x"BB",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B2",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FA",x"D5",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"FF",x"F5",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"BB",x"13",
x"13",x"57",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B1",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D5",x"D1",
x"D1",x"D1",x"FF",x"F6",x"FF",x"D1",x"D1",x"FB",x"FA",x"D1",x"FF",x"FF",x"FF",x"9B",x"13",x"13",
x"13",x"13",x"9B",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AD",x"44",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FA",x"FA",x"FF",x"FA",x"FF",x"F5",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"77",x"13",x"13",x"13",
x"13",x"13",x"37",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FB",x"FF",x"9B",x"57",x"9B",x"DF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"F6",x"FF",x"F6",x"D1",x"F6",x"FF",x"FF",x"FF",x"57",x"13",x"13",x"13",x"13",
x"13",x"13",x"13",x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"DF",x"13",x"13",x"13",x"13",x"13",x"33",
x"77",x"FF",x"FF",x"D1",x"F6",x"D5",x"D1",x"D1",x"FA",x"FB",x"FF",x"33",x"13",x"13",x"13",x"13",
x"13",x"13",x"13",x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"77",x"13",x"13",x"13",x"13",x"13",x"13",
x"13",x"BF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"57",x"13",x"13",x"13",x"13",
x"13",x"13",x"57",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"91",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"37",x"13",x"13",x"13",x"13",x"13",x"13",
x"13",x"9B",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"BB",x"13",x"13",x"13",x"13",
x"13",x"13",x"DF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"57",x"13",x"13",x"13",x"13",x"13",x"13",
x"13",x"BB",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"77",x"13",x"13",x"13",
x"13",x"BB",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B1",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"9B",x"13",x"13",x"13",x"13",x"13",x"13",
x"13",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"DF",x"9B",x"9B",
x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B6",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",x"44",x"68",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C8",x"CC",x"D1",x"D1",x"FF",x"FF",x"33",x"13",x"13",x"13",x"13",x"13",
x"77",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",
x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"D6",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"64",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C0",x"C4",x"D1",x"D1",x"FA",x"FF",x"DF",x"33",x"13",x"13",x"13",x"77",
x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"FB",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"44",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C0",x"C0",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"BB",x"9B",x"DF",x"FF",
x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"68",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"88",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C0",x"C0",x"CC",x"D1",x"D1",x"D1",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"8D",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"68",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C4",x"C0",x"C4",x"D1",x"D1",x"D1",x"D1",x"D5",x"FA",x"FA",x"FA",x"D5",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"B2",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"64",x"B1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"CD",x"C0",x"C0",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"FB",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"88",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",x"C0",x"C0",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"68",x"FF",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"64",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",x"C0",x"C0",x"C4",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"B2",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"44",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C4",x"C0",x"C0",x"C0",x"C4",x"C8",x"CC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CD",x"CC",x"CD",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"68",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C4",x"C0",x"C0",x"C0",x"C0",x"C0",
x"C0",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C0",x"C0",x"C0",x"C0",x"C8",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"8D",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"44",
x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C8",x"C4",x"C4",
x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C4",x"C8",x"C8",x"CD",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",
x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"CD",x"CD",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",
x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",
x"64",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"B1",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"68",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"89",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"DA",x"B1",x"8D",x"8D",x"B2",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FF",x"68",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"68",x"64",x"44",x"44",x"44",x"44",x"64",x"B1",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"DB",x"64",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"88",x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"B1",x"64",x"44",x"68",x"B2",x"D6",x"D6",x"B1",x"64",x"44",x"8D",x"FF",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"DB",x"64",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"B1",x"44",x"64",x"D6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"89",x"44",x"8D",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"DB",x"68",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"64",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"D6",x"44",x"64",x"C0",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"68",x"44",
x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"B2",x"64",x"64",x"44",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",
x"64",x"64",x"64",x"8D",x"DB",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FF",x"68",x"64",x"C0",x"C0",x"C9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"64",
x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FB",x"89",x"44",x"64",x"AC",x"88",x"64",x"44",x"64",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",
x"88",x"D1",x"D1",x"88",x"64",x"B1",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"B2",x"44",x"A4",x"C0",x"C0",x"C0",x"ED",x"FB",x"D6",x"FF",x"FF",x"FB",x"F6",x"ED",x"84",
x"44",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"D6",x"64",x"44",x"68",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"AD",
x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"68",x"B6",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"68",x"68",x"C4",x"C0",x"C0",x"C0",x"84",x"64",x"44",x"64",x"A9",x"C0",x"C0",x"C0",x"C0",
x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",
x"8D",x"64",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"8D",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"DA",x"44",x"B2",x"F6",x"C0",x"C0",x"84",x"44",x"68",x"8D",x"64",x"64",x"C0",x"C0",x"C0",x"C0",
x"84",x"44",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"89",
x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"64",x"64",x"B2",x"FF",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"B1",x"64",x"DB",x"FF",x"F2",x"A0",x"64",x"68",x"FF",x"FF",x"D6",x"44",x"84",x"C0",x"C0",x"C0",
x"A0",x"64",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"68",x"44",
x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"8D",x"68",x"FF",x"FF",x"FF",x"B1",x"44",x"D6",x"E0",x"E0",x"FF",x"8D",x"64",x"C9",x"F6",x"FB",
x"FB",x"68",x"68",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"64",x"44",x"64",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FA",x"FA",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"64",x"D6",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"68",x"89",x"FF",x"FF",x"FF",x"8D",x"64",x"FF",x"E0",x"E0",x"E0",x"D6",x"44",x"B2",x"FF",x"FF",
x"FF",x"8D",x"64",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"B6",x"64",x"44",x"68",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",
x"D1",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"64",x"64",x"B2",x"FF",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"64",x"8D",x"FF",x"FF",x"FF",x"8D",x"68",x"FF",x"E0",x"E0",x"E0",x"FF",x"64",x"68",x"FF",x"FF",
x"FF",x"D6",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"B2",x"64",x"44",x"68",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"B1",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"64",x"8D",x"FF",x"FF",x"FF",x"8D",x"64",x"FF",x"E0",x"E0",x"FF",x"FF",x"8D",x"64",x"FF",x"FF",
x"FF",x"FB",x"64",x"B1",x"E0",x"E0",x"E0",x"E0",x"FF",x"B1",x"44",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",
x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"68",x"89",x"FF",x"FF",x"FF",x"D6",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"D6",x"FF",
x"FF",x"FF",x"68",x"68",x"E0",x"E0",x"E0",x"FF",x"8D",x"44",x"64",x"8C",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FB",x"FF",x"FA",x"FA",x"FF",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"B1",x"64",
x"64",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"8D",x"68",x"FF",x"FF",x"FF",x"FB",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"8D",x"FF",
x"FF",x"FF",x"8D",x"64",x"FF",x"E0",x"FF",x"8D",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"D1",x"FF",x"F5",x"F6",x"FF",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",
x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"B2",x"44",x"A4",x"C9",x"C4",x"C4",x"64",x"64",x"FF",x"E0",x"E0",x"E0",x"FF",x"68",x"68",x"FF",
x"FF",x"FF",x"B6",x"44",x"DA",x"FF",x"89",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FA",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"68",x"64",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"DB",x"64",x"84",x"C0",x"C0",x"C0",x"84",x"44",x"FB",x"E0",x"E0",x"E0",x"E0",x"91",x"64",x"FF",
x"FF",x"FF",x"FB",x"44",x"8D",x"68",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FB",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"64",x"D1",x"D1",x"AC",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"8C",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"68",x"64",x"A0",x"C0",x"C0",x"84",x"44",x"FF",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"A4",
x"C4",x"C9",x"F2",x"64",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FB",x"FB",x"FA",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"AC",x"AC",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"DA",x"64",x"64",x"A4",x"84",x"64",x"68",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"84",
x"C0",x"C0",x"C0",x"64",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"64",x"88",x"64",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FF",x"B1",x"64",x"44",x"44",x"64",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"64",
x"C0",x"C0",x"C0",x"84",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"68",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"D6",x"91",x"B2",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"64",
x"C4",x"C0",x"C0",x"A0",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"68",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"D5",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"88",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"44",
x"D6",x"FF",x"FB",x"F2",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"8C",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",x"44",
x"B2",x"FF",x"FF",x"FF",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"8C",x"44",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"8D",x"44",
x"8D",x"FF",x"FF",x"FF",x"B1",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"68",x"44",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"64",x"44",
x"68",x"FF",x"FF",x"FF",x"D6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"B1",x"64",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"64",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"64",
x"64",x"FF",x"FF",x"FF",x"FB",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"F5",x"FF",x"D1",x"FA",x"FF",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",
x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"64",x"68",x"AC",
x"44",x"D6",x"FF",x"FF",x"FF",x"68",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"44",x"68",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FA",x"F5",x"FF",x"FA",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",
x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",
x"44",x"B1",x"FF",x"FF",x"FF",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"68",x"44",x"64",x"B1",x"FF",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",
x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"64",x"D1",x"D1",
x"64",x"89",x"FF",x"FF",x"FF",x"B2",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",
x"64",x"44",x"68",x"D6",x"E0",x"FB",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",
x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"88",x"D1",x"D1",
x"88",x"64",x"FF",x"FF",x"FF",x"DB",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"44",
x"44",x"8D",x"FF",x"E0",x"E0",x"D6",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"F6",x"D5",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"68",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"AC",x"D1",x"D1",
x"8C",x"44",x"C9",x"E9",x"F2",x"F6",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"44",x"64",
x"B6",x"FF",x"E0",x"E0",x"E0",x"B2",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"64",x"DB",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"AC",x"D1",x"D1",
x"AC",x"44",x"A4",x"C0",x"C0",x"C0",x"64",x"64",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"8D",x"FB",
x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"68",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"64",x"B6",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"AC",x"D1",x"D1",
x"D1",x"64",x"84",x"C0",x"C0",x"C0",x"84",x"44",x"AC",x"68",x"64",x"44",x"68",x"D6",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"68",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"AC",x"AC",x"8C",x"64",x"44",x"44",x"B2",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",x"44",x"68",x"D1",x"D1",
x"D1",x"68",x"64",x"C0",x"C0",x"C0",x"A4",x"44",x"44",x"44",x"64",x"B1",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"44",x"44",x"64",x"B6",x"FF",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"44",x"68",x"AC",
x"D1",x"88",x"64",x"CD",x"C9",x"C4",x"C0",x"64",x"64",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"FB",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"64",x"64",x"64",x"8D",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"64",x"44",x"44",
x"44",x"44",x"44",x"D6",x"FF",x"FF",x"F6",x"68",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"DA",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",x"D6",x"FB",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"8D",x"64",
x"64",x"64",x"44",x"B2",x"FF",x"FF",x"FF",x"8D",x"64",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"B6",x"44",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",
x"FB",x"DB",x"64",x"8D",x"FF",x"FF",x"FF",x"B6",x"44",x"DA",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"91",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"8D",x"64",x"FF",x"FF",x"FF",x"DB",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B2",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"B1",x"44",x"FB",x"FF",x"FF",x"FF",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"68",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"B1",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"D6",x"44",x"B6",x"FF",x"FF",x"FF",x"8D",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"64",x"8D",x"FF",x"FF",x"FF",x"B2",x"44",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FB",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"68",x"68",x"FF",x"FF",x"FF",x"DA",x"44",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"DA",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"8D",x"64",x"FF",x"FF",x"FF",x"FF",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"B6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"68",x"68",x"88",x"8C",x"AD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"B6",x"44",x"D6",x"FF",x"FF",x"FF",x"68",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"B1",x"44",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"44",x"44",x"44",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FB",x"44",x"89",x"F2",x"FB",x"FF",x"B1",x"64",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"64",x"B6",x"D6",x"D6",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"64",x"64",x"C0",x"C0",x"C9",x"AD",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"88",x"68",x"FF",x"E0",x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"8D",x"64",x"C0",x"C0",x"C0",x"C0",x"64",x"B1",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"68",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"64",x"B1",x"E0",x"E0",x"E0",x"8D",x"44",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"89",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"A0",x"C0",x"C0",x"C0",x"64",x"68",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"DB",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"89",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"DA",x"44",x"A8",x"C9",x"C0",x"C0",x"84",x"64",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"DB",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"68",x"FF",x"E0",x"E0",x"E0",x"91",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"89",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"8D",x"FF",x"FF",x"F2",x"A4",x"44",x"DA",x"E0",x"E0",x"E0",
x"E0",x"E0",x"D6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"89",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"68",x"68",x"FF",x"FF",x"FF",x"DB",x"44",x"B2",x"E0",x"E0",x"E0",
x"E0",x"E0",x"B2",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"89",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"B1",x"64",x"FB",x"FF",x"FF",x"FF",x"64",x"8D",x"E0",x"E0",x"E0",
x"E0",x"E0",x"8D",x"44",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"88",x"64",x"FF",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"D6",x"FF",x"FF",x"FF",x"8D",x"68",x"FF",x"E0",x"E0",
x"E0",x"E0",x"8D",x"44",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"B1",x"FF",x"FF",x"FF",x"B1",x"44",x"FB",x"E0",x"E0",
x"E0",x"FF",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"64",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"68",x"FF",x"FF",x"FF",x"D6",x"44",x"B6",x"E0",x"E0",
x"E0",x"FF",x"64",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"88",x"64",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"64",x"FF",x"FF",x"FF",x"FF",x"44",x"8D",x"E0",x"E0",
x"E0",x"FB",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B2",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"DB",x"FF",x"FF",x"FF",x"68",x"68",x"FF",x"E0",
x"E0",x"D6",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FB",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",x"44",x"B6",x"FF",x"FF",x"FF",x"8D",x"64",x"FF",x"E0",
x"E0",x"B6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",
x"44",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"8D",x"FB",x"FF",x"FF",x"B6",x"44",x"DB",x"E0",
x"E0",x"B1",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",
x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"64",x"C0",x"C4",x"ED",x"CD",x"44",x"D6",x"E0",
x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",
x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"91",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"91",x"64",x"C0",x"C0",x"C0",x"A0",x"44",x"B6",x"E0",
x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",
x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"84",x"C0",x"C0",x"A0",x"44",x"B6",x"E0",
x"E0",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"44",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"64",x"A0",x"C0",x"84",x"44",x"DB",x"E0",
x"E0",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"64",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"64",x"64",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"44",x"64",x"64",x"44",x"68",x"FF",x"E0",
x"E0",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",x"B6",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"64",x"AD",x"D1",x"D1",
x"D1",x"8C",x"64",x"44",x"B2",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"B2",x"64",x"44",x"68",x"FF",x"E0",x"E0",
x"E0",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"FF",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"44",x"64",x"68",x"88",
x"64",x"44",x"44",x"B1",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",
x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"8D",x"64",x"44",x"44",
x"44",x"64",x"B6",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"91",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"DB",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"B2",x"B1",
x"D6",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"D6",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"8D",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FF",x"64",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"FB",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"B1",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"64",x"D6",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"68",x"44",x"64",x"88",x"88",x"68",x"64",x"64",x"B6",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FB",x"68",x"44",x"44",x"44",x"44",x"68",x"DA",x"FF",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"FF",x"B6",x"8D",x"8D",x"D6",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0");
  
	constant cookieL : characterImage := (
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"40",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"64",
x"64",x"68",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"68",x"64",x"64",x"44",x"44",
x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"88",x"AC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"88",
x"68",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"64",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"88",x"68",x"64",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"64",x"88",x"D0",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"F6",x"F6",x"F6",x"F6",x"F6",x"F5",x"F5",
x"F5",x"F5",x"D1",x"D1",x"AC",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"D6",x"91",x"8D",x"DB",x"FF",x"B6",x"24",x"24",x"24",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"40",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DB",
x"92",x"92",x"49",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"92",x"24",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D5",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FA",x"F5",x"F6",x"FA",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"24",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"FF",x"FF",x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"B1",x"8D",x"DA",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"24",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",
x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"F5",x"FB",x"FF",x"FF",x"FF",x"FF",x"FB",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"6D",
x"49",x"DB",x"FF",x"FF",x"FF",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"F5",x"D1",x"D1",
x"D1",x"D1",x"F5",x"FB",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",
x"F5",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"8D",x"D5",
x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FA",x"FA",x"F5",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"88",
x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"6D",x"92",x"FF",x"FF",x"FF",x"FF",x"FF",x"F2",x"60",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"64",x"D6",x"FF",
x"FF",x"FF",x"FF",x"FA",x"F6",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FA",x"F6",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",
x"64",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F2",x"C4",x"C4",x"A0",x"20",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"FA",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FA",x"D1",x"F5",x"F6",x"FB",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",
x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"49",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F2",x"C4",x"C4",x"C4",x"C4",x"80",x"40",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"44",x"AC",x"D1",x"D1",
x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"F6",x"F5",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"F5",x"FA",
x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",
x"D1",x"68",x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"FB",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"ED",x"C4",x"C4",x"C4",x"C4",x"C4",x"CD",x"6D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",
x"F6",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F5",x"F6",x"FA",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",
x"D1",x"AC",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"80",x"C4",x"F2",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"ED",x"C4",x"C4",x"C4",x"C4",x"C4",x"F6",x"FF",x"49",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FA",x"F5",x"F5",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"F5",x"F5",x"F5",x"F5",x"F5",x"D1",x"D1",x"D1",
x"D1",x"D1",x"64",x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"C4",x"C4",x"C4",x"C9",
x"F6",x"FF",x"FF",x"FF",x"DB",x"DB",x"DB",x"CD",x"C4",x"C4",x"C4",x"C4",x"C4",x"FB",x"FF",x"FF",
x"49",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"60",x"C4",x"C4",x"C4",x"C4",
x"C4",x"ED",x"B2",x"49",x"E0",x"E0",x"E0",x"20",x"80",x"C4",x"C4",x"C4",x"C9",x"FF",x"FF",x"FF",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D0",x"64",x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"C4",x"C4",x"C4",x"C4",x"C4",
x"C4",x"80",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"A4",x"C4",x"ED",x"FF",x"FF",x"FF",
x"FF",x"6D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",x"FA",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"C4",x"C4",x"C4",x"C4",x"C4",
x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"C4",x"F6",x"FF",x"FF",x"FF",
x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FB",x"D1",x"FA",x"F5",x"F6",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"FB",x"F2",x"C9",x"C4",x"C4",
x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"A9",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"D1",x"FA",x"F5",x"D1",
x"FF",x"F5",x"F5",x"FA",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"F5",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"40",x"E0",x"E0",x"E0",x"24",x"FF",x"FF",x"FB",x"ED",x"C4",
x"A4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"6D",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"D1",x"FA",x"F5",x"F5",
x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"F5",x"F5",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"F5",x"FA",x"FB",x"FF",x"FF",x"FB",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"24",x"FF",x"FF",x"FF",x"FF",x"FB",
x"ED",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"D1",x"FF",x"F6",x"F5",
x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",
x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"E0",x"E0",x"E0",x"24",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"FF",x"FF",x"FF",
x"FF",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"CC",x"D1",x"D1",x"F5",x"FB",x"FB",
x"F6",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"D1",x"FF",x"F6",x"F6",
x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"20",x"E0",x"E0",x"24",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"6D",x"FF",x"FF",x"FF",
x"FF",x"FF",x"92",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",
x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"D1",x"FF",x"F6",x"FA",
x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D0",x"64",x"44",x"20",x"E0",x"E0",x"24",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"92",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",
x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"F5",x"D1",x"D1",x"F6",x"FF",x"FF",x"D1",x"FF",x"F6",x"FA",
x"FF",x"FA",x"D1",x"D1",x"F5",x"F5",x"F6",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"DB",x"FF",x"FF",x"FF",x"FF",
x"FF",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FF",
x"B6",x"49",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"F5",x"FA",x"FF",x"FF",x"D1",x"FF",x"F6",x"F6",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"92",x"FF",x"FF",x"FF",x"FF",
x"F2",x"A9",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"49",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"F5",x"FF",x"F5",x"F5",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"BB",x"9B",x"FF",x"FF",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"92",x"FF",x"FF",x"FF",x"ED",
x"C4",x"C4",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",
x"FF",x"DF",x"77",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"FA",x"D1",x"D1",
x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"BB",x"97",x"57",x"33",x"12",x"12",x"FF",x"FF",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"E9",x"C4",
x"C4",x"C4",x"60",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",
x"FF",x"9B",x"0E",x"12",x"53",x"9B",x"BB",x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"FB",x"FF",x"DF",x"33",x"12",x"0E",x"0E",x"0E",x"0E",x"0E",x"33",x"FF",x"FF",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"92",x"ED",x"C4",x"C4",
x"C4",x"C4",x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",
x"FF",x"9B",x"0E",x"0E",x"0E",x"0E",x"12",x"DF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"FA",x"FF",x"FF",x"33",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"77",x"FF",x"FA",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"40",x"C4",x"C4",x"C4",
x"C4",x"C4",x"C4",x"92",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",
x"FF",x"BB",x"0E",x"0E",x"0E",x"0E",x"33",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F6",x"FF",x"FF",x"57",x"0E",x"0E",x"0E",x"0E",x"0E",x"12",x"BB",x"FF",x"F6",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"C4",x"C4",x"C4",
x"C4",x"C9",x"FB",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"CC",x"D1",x"D1",x"D1",x"D1",x"F5",
x"FF",x"DB",x"0E",x"0E",x"0E",x"0E",x"9B",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F5",x"FF",x"FF",x"9B",x"0E",x"0E",x"0E",x"0E",x"0E",x"33",x"FF",x"FF",x"F5",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"80",x"C4",x"C4",
x"C9",x"FB",x"FF",x"FF",x"24",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"F5",
x"FF",x"FF",x"33",x"0E",x"0E",x"12",x"DF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"33",x"0E",x"0E",x"0E",x"0E",x"9B",x"FF",x"FF",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"C4",x"C9",
x"FB",x"FF",x"FF",x"FF",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"FB",x"FF",x"BB",x"33",x"33",x"77",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"BB",x"33",x"12",x"12",x"77",x"FF",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"A4",x"F6",
x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",
x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"DF",x"BB",x"BB",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"69",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"49",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",
x"FF",x"FF",x"FF",x"FF",x"FF",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F5",x"F6",x"F6",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FA",x"FB",x"FB",x"FA",x"F5",x"CD",x"CC",x"C8",x"C8",
x"C8",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CD",x"C8",x"C4",x"C4",x"C4",x"C4",x"C4",
x"C4",x"C4",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"92",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"6D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C8",x"C8",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",
x"C4",x"C4",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"CC",x"C8",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C8",x"CC",x"D1",x"C8",
x"C4",x"C4",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"CC",x"64",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"92",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"69",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CD",x"C8",x"C8",x"C4",
x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C8",x"CC",x"CD",x"D1",x"D1",x"D1",x"D1",x"C8",
x"C4",x"C4",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"68",x"DA",x"FF",x"FF",x"FF",x"F2",x"C4",x"64",x"44",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C8",x"C4",x"C4",x"C4",x"C4",x"C4",
x"C4",x"C4",x"C4",x"C8",x"C8",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",
x"C4",x"C4",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"64",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",
x"44",x"8D",x"FF",x"FF",x"F2",x"C4",x"C4",x"84",x"44",x"44",x"44",x"44",x"20",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CD",x"C4",x"C4",x"C4",x"C4",x"C4",x"C8",x"C8",
x"CC",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",
x"C4",x"C4",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"44",x"44",x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"44",x"44",x"44",x"44",
x"64",x"88",x"DB",x"F2",x"C4",x"C4",x"C4",x"C4",x"88",x"68",x"44",x"44",x"44",x"20",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C4",x"C4",x"C4",x"C4",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",
x"C4",x"C4",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"CC",x"64",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"64",x"88",x"AC",
x"D1",x"D1",x"F1",x"C4",x"C4",x"C4",x"C4",x"C4",x"CD",x"D1",x"88",x"44",x"44",x"44",x"20",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"8C",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C4",x"C4",x"C4",x"C8",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C4",
x"C4",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"88",x"44",x"44",x"44",x"44",x"E0",x"20",x"44",x"44",x"44",x"64",x"68",x"8C",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"C4",x"C4",x"C4",x"C4",x"ED",x"FA",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",x"C4",x"C4",x"C4",x"CC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C4",
x"C4",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",
x"44",x"44",x"44",x"44",x"20",x"44",x"44",x"44",x"44",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"C8",x"C4",x"C4",x"ED",x"FF",x"FF",x"F5",x"D1",x"D1",x"64",x"44",x"44",x"20",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",x"C4",x"C4",x"C4",x"CC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CD",x"C4",
x"C4",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",
x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"CC",x"C4",x"C9",x"FB",x"FF",x"FF",x"FA",x"D1",x"D1",x"88",x"44",x"44",x"20",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"44",
x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C4",x"C4",x"C4",x"C4",
x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",x"C4",
x"C4",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",
x"44",x"44",x"44",x"44",x"44",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C8",x"F6",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"AC",x"44",x"44",x"20",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",x"C4",x"C4",
x"C4",x"C4",x"C8",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C4",x"C4",
x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",
x"44",x"44",x"44",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"F1",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"AC",x"44",x"44",x"20",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",
x"44",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C4",
x"C4",x"C4",x"C4",x"C4",x"C4",x"C8",x"C8",x"CC",x"CC",x"CC",x"CC",x"CC",x"C8",x"C4",x"C4",x"C8",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",
x"44",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"88",x"44",x"44",x"20",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"C8",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C8",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"64",x"88",
x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"68",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"44",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"CD",x"C8",x"C8",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"CC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"64",x"8C",x"AC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"D6",x"44",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"20",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"20",x"E0",x"20",x"44",x"44",x"88",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"CD",x"CC",x"CC",x"CC",x"CC",x"CC",x"CD",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"DB",x"64",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"69",x"44",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"44",x"64",x"68",x"88",x"AC",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D0",x"AC",x"AC",x"88",
x"88",x"68",x"64",x"44",x"44",x"44",x"44",x"44",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"D6",x"20",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",
x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"AC",x"88",x"68",x"64",x"64",x"64",x"68",x"8C",x"D0",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"ED",x"40",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"44",x"88",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"AC",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"F2",x"C4",x"A0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"68",x"FF",x"FF",x"FB",x"C4",x"C4",x"C4",x"40",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"AC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"D6",x"FF",x"C9",x"C4",x"C4",x"C4",x"60",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"CC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D0",x"88",x"64",x"44",x"44",x"44",x"8D",x"F2",x"C4",x"C4",x"C4",x"C4",x"C4",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"64",x"44",x"44",x"44",x"44",x"E0",x"40",x"C4",x"C4",x"C4",x"C4",x"C4",x"F6",x"49",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",
x"68",x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"80",x"C4",x"C4",x"C4",x"F2",x"FF",x"B6",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"AC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"88",x"44",
x"44",x"44",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"60",x"C4",x"C4",x"C9",x"FF",x"FF",x"FF",
x"49",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"44",x"8C",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"D1",x"F5",x"FF",x"FA",x"D1",x"F6",x"FF",x"F6",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"88",x"64",x"44",x"44",
x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C4",x"C4",x"F6",x"FF",x"FF",x"FF",
x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"F5",x"F5",x"FF",x"FF",x"F5",x"FA",x"FF",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"44",x"44",x"44",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"80",x"ED",x"FF",x"FF",x"FF",x"FF",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"44",x"88",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"44",x"44",x"44",x"44",x"44",x"20",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"49",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"92",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",
x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"44",x"44",x"44",x"44",x"20",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FF",x"FF",x"FF",x"FF",
x"FF",x"92",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"44",
x"44",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FB",x"FB",x"F6",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"64",x"44",x"44",x"44",x"44",x"40",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"92",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",
x"44",x"44",x"64",x"88",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"F5",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"88",x"64",x"44",x"44",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"92",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"44",x"44",x"44",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"68",x"44",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"40",x"44",x"44",x"44",x"44",x"44",x"64",x"88",x"AC",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"6D",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"6D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"20",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"88",x"88",x"AC",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FB",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FF",x"FF",
x"FF",x"FF",x"FF",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"64",
x"64",x"64",x"68",x"88",x"88",x"AC",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"CC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FF",x"FF",
x"FF",x"FF",x"F6",x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"E0",x"40",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"88",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"24",x"FF",x"FF",
x"FF",x"F6",x"C4",x"C4",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"24",x"FF",x"FF",
x"FB",x"C9",x"C4",x"C4",x"80",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"92",x"FF",
x"ED",x"C4",x"C4",x"C4",x"C4",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"F5",x"F5",x"FF",x"FF",x"F5",x"F5",x"FF",
x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"92",x"ED",
x"C4",x"C4",x"C4",x"C4",x"C9",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"F6",x"F5",x"FF",x"FF",x"F5",x"F6",x"FF",
x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"A0",
x"C4",x"C4",x"C4",x"C4",x"FB",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",
x"C4",x"C4",x"C4",x"F6",x"FF",x"FF",x"92",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"40",x"40",x"44",x"44",x"88",x"AC",x"AC",x"AC",
x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"A0",x"C4",x"ED",x"FF",x"FF",x"FF",x"92",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"64",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FA",x"FA",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"80",x"C9",x"FB",x"FF",x"FF",x"FF",x"FF",x"24",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"40",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"64",x"64",x"64",x"64",x"68",
x"88",x"8C",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"F5",x"F5",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"92",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"44",x"44",x"44",x"64",x"88",x"8C",x"AC",x"AC",x"AC",x"AC",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"DB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"44",x"88",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"6D",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"92",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",
x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"20",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"49",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",
x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"DB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",
x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",
x"44",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"8C",x"88",x"88",x"68",x"68",x"64",x"64",x"64",x"64",
x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"20",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"92",x"FF",x"FF",x"FF",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"6D",x"FF",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"40",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"44",x"44",x"44",x"44",x"40",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"40",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"44",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D0",x"64",x"44",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"40",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"20",x"44",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",
x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",
x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"44",x"64",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",
x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",
x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"44",x"68",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"88",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"44",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"44",x"68",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"8C",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"88",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",
x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"88",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"64",
x"88",x"8C",x"8C",x"8C",x"88",x"44",x"44",x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",
x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",
x"44",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"44",x"44",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"40",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"8C",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"8C",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"40",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"20",x"44",x"44",x"64",x"88",x"AC",x"AC",x"AC",x"AC",x"88",
x"64",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0");
	
		constant cookieR : characterImage := (
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"44",x"44",x"44",x"64",x"64",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"64",
x"64",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"64",x"68",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"CC",x"AC",x"88",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"88",
x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"64",x"88",x"AC",x"D1",x"D1",
x"D1",x"D5",x"F5",x"F5",x"F5",x"F5",x"F5",x"F5",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"88",x"64",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"BB",x"DB",x"92",x"E0",x"8D",x"B2",x"FA",x"FA",x"FA",x"FB",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"F1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"72",
x"96",x"96",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"96",x"DB",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FA",x"FB",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FB",x"B6",x"D6",x"F6",x"F5",x"F5",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",x"FA",x"FF",x"FF",
x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",
x"DB",x"BA",x"B6",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",
x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"71",x"E0",x"E0",
x"E0",x"E0",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",
x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"68",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"44",x"64",x"CC",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",
x"D1",x"F5",x"F6",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"64",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"AD",x"DB",x"DB",x"DB",x"DB",x"DB",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"88",x"D1",x"D1",x"D1",x"F5",x"FB",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"F5",x"FA",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"64",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"84",x"C4",x"C4",x"F2",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"92",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"68",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"F5",x"FA",x"FA",
x"FF",x"FF",x"D6",x"64",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"A4",x"C4",x"C4",x"C4",x"F2",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",
x"44",x"AC",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"F5",x"F5",x"FA",x"FF",x"FF",x"FB",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FA",x"FB",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"D5",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"A9",x"C4",x"C4",x"C4",x"C4",x"C4",x"ED",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",
x"68",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",x"F5",x"FB",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FA",x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"DB",x"F6",x"C4",x"C4",x"C4",x"C4",x"C4",x"ED",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FB",x"ED",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"64",
x"AC",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FA",x"F6",
x"F5",x"D1",x"D1",x"D1",x"D1",x"F5",x"FB",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"F5",x"FA",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"F6",
x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"DB",x"FF",x"FB",x"C4",x"C4",x"C4",x"C4",x"C4",x"ED",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"F2",x"C4",x"C4",x"A4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",
x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",x"FA",x"FA",x"FA",x"FA",x"F6",x"F5",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"F5",x"F6",x"FA",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"BA",x"FF",x"FF",x"FF",x"C9",x"C4",x"C4",x"C4",x"C4",x"A9",x"E0",x"E0",x"E0",x"DB",x"FF",
x"F6",x"C9",x"C4",x"C4",x"C4",x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"8C",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FA",x"D5",x"F5",x"FA",x"FB",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"F6",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"CC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FF",x"FF",x"FF",x"FF",x"ED",x"C4",x"C4",x"A4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"A4",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"96",x"FF",x"FF",x"FF",x"FF",x"F6",x"C4",x"88",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"C9",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"C4",x"C4",x"C4",x"C4",x"C9",x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"64",x"AC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FA",x"FB",x"F5",x"F6",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"C4",x"C4",x"C4",x"F2",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"68",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FA",
x"FF",x"F5",x"D1",x"FA",x"D1",x"FA",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"72",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"A4",x"ED",x"FB",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"8C",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FB",x"FA",x"F5",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FA",x"FA",x"FA",x"FA",x"FA",x"F6",x"F5",x"D1",x"D1",x"D1",
x"FF",x"F6",x"D5",x"FB",x"D1",x"FA",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"BA",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"44",x"64",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",
x"FF",x"FA",x"F5",x"FF",x"D1",x"FA",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"BA",
x"FF",x"FF",x"FF",x"FF",x"FF",x"BA",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D0",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FA",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",
x"FF",x"FA",x"F5",x"FF",x"D1",x"FA",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"F5",x"F5",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"71",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",
x"FF",x"FA",x"F5",x"FF",x"D1",x"FB",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",
x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"CC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"DB",x"FF",x"FF",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FB",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",
x"FF",x"FB",x"F5",x"FF",x"F5",x"FB",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"F6",x"FA",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"DF",x"BA",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"D6",x"FB",x"FF",x"FF",x"FF",x"FF",x"B6",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FA",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FA",x"F6",x"F6",x"FB",
x"FF",x"FB",x"F5",x"FF",x"F5",x"FB",x"FF",x"FA",x"D1",x"F5",x"F6",x"FB",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"A4",x"C9",x"FB",x"FF",x"FF",x"FF",x"96",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"F5",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FA",x"F5",x"FF",x"F5",x"FA",x"FF",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"68",
x"C4",x"C4",x"C9",x"F6",x"FF",x"FF",x"96",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F6",x"FF",x"97",x"57",x"9B",x"BB",x"DF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"F5",x"D1",x"FA",x"F5",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DF",x"FF",
x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"A4",
x"C4",x"C4",x"C4",x"C4",x"FB",x"DF",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F6",x"FF",x"77",x"0E",x"0E",x"0E",x"33",x"57",x"77",x"9B",x"DF",x"FF",x"FF",x"FA",
x"D1",x"D1",x"D1",x"F5",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"DB",x"77",x"33",x"9B",
x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C4",
x"C4",x"C4",x"C4",x"C4",x"C9",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F5",x"FF",x"BB",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"0E",x"9B",x"FF",x"FF",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"77",x"33",x"12",x"0E",x"0E",x"9B",
x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"BA",x"ED",
x"C4",x"C4",x"C4",x"C4",x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F5",x"FF",x"DF",x"12",x"0E",x"0E",x"0E",x"0E",x"0E",x"12",x"DB",x"FF",x"FF",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"33",x"0E",x"0E",x"0E",x"0E",x"9B",
x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FF",
x"ED",x"C4",x"C4",x"C4",x"A4",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"FF",x"FF",x"53",x"0E",x"0E",x"0E",x"0E",x"0E",x"33",x"FF",x"FF",x"FA",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"77",x"0E",x"0E",x"0E",x"0E",x"9B",
x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"CC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"72",x"FF",x"FF",
x"FF",x"ED",x"C4",x"C4",x"88",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"FA",x"FF",x"9B",x"12",x"0E",x"0E",x"0E",x"0E",x"77",x"FF",x"FF",x"F6",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"DB",x"12",x"0E",x"0E",x"12",x"BB",
x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",
x"FF",x"FF",x"C9",x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"57",x"0E",x"0E",x"0E",x"33",x"DF",x"FF",x"FF",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"57",x"0E",x"0E",x"57",x"FF",
x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FB",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"DF",x"77",x"33",x"53",x"BB",x"FF",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"BB",x"77",x"77",x"DF",x"FF",
x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"88",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FB",x"F5",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"68",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CD",
x"C4",x"C4",x"C4",x"C4",x"C8",x"CC",x"D1",x"F6",x"F6",x"F6",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"72",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",
x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C8",x"CC",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"DF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"88",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",
x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C8",x"C8",x"CC",x"CD",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D1",x"FF",x"FF",x"FF",x"FF",
x"FF",x"96",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",
x"C4",x"C4",x"CD",x"D1",x"CC",x"C8",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C8",
x"C8",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"64",x"C4",x"ED",x"FF",x"FF",x"FF",
x"B2",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",
x"C4",x"C4",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C8",x"C8",x"C4",x"C4",x"C4",x"C4",x"C4",
x"C4",x"C4",x"C4",x"C4",x"C8",x"CC",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"84",x"C4",x"C4",x"ED",x"FF",x"FF",
x"68",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"68",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",
x"C4",x"C4",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C8",x"C8",x"C4",
x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C8",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"88",x"AC",x"C4",x"C4",x"C4",x"C4",x"ED",x"DA",
x"8C",x"68",x"64",x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",
x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",
x"C4",x"C4",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"CD",x"CC",x"C8",x"C4",x"C4",x"C4",x"C4",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"8C",x"D1",x"D1",x"C4",x"C4",x"C4",x"C4",x"C4",x"D1",
x"D1",x"D1",x"AC",x"88",x"64",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",
x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",
x"C4",x"C4",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C8",x"C4",x"C4",x"C4",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"68",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"44",x"8C",x"D1",x"D1",x"FA",x"F2",x"C4",x"C4",x"C4",x"C4",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"88",x"64",x"44",x"44",x"44",x"E0",x"E0",x"44",x"44",x"44",
x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CD",
x"C4",x"C4",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"C8",x"C4",x"C4",x"C4",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"F5",x"FF",x"FF",x"ED",x"C4",x"C4",x"C8",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"88",x"44",x"44",x"44",x"44",x"48",x"44",x"44",
x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"C4",x"C4",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"CC",x"C4",x"C4",x"C4",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"ED",x"C4",x"CD",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D0",x"88",x"64",x"44",x"44",x"44",x"44",
x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"C8",x"C4",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"CC",x"C4",x"C4",x"C4",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"8C",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FB",x"C9",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"44",x"44",x"44",
x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"CC",x"C4",x"C4",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"C8",x"C4",x"C4",x"C4",x"C4",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"8C",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"44",
x"44",x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"C8",x"C4",x"C4",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CD",x"C8",x"C4",
x"C4",x"C4",x"C4",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",
x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",
x"68",x"44",x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"CD",x"C4",x"C4",x"C4",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C4",x"C4",x"C4",x"C4",
x"C4",x"C4",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",
x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"88",x"64",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"CD",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",
x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"44",x"B1",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"88",x"64",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"CD",x"C8",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C8",x"C8",x"CD",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"44",x"64",x"D6",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"88",x"D0",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CD",x"CC",x"CC",x"CC",x"CC",x"CD",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"88",x"44",x"44",x"44",x"E0",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"44",x"68",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"44",x"44",x"44",x"44",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"88",x"44",x"44",x"44",x"44",x"44",x"64",x"68",
x"88",x"8C",x"AC",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D0",x"AC",x"88",x"68",x"44",
x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"64",x"64",x"68",x"68",x"88",x"AC",x"CC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",
x"64",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"A4",x"C4",x"ED",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"AC",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"C4",x"C4",x"C4",x"F6",x"FF",x"FF",x"68",x"68",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"C4",x"C4",x"C4",x"C9",x"FF",x"D6",x"44",x"44",x"64",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FB",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"A4",x"C4",x"C4",x"C4",x"C4",x"F2",x"8D",x"44",x"44",x"44",x"64",x"88",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FB",x"C9",x"C4",x"C4",x"C4",x"C4",x"E0",x"E0",x"44",x"44",x"44",x"44",x"64",
x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"BA",x"FF",x"F2",x"C4",x"C4",x"C4",x"A4",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",
x"44",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"FF",x"FF",x"C9",x"C4",x"C4",x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"44",x"44",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"BA",x"FF",x"FF",x"FF",x"F6",x"C4",x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",
x"44",x"44",x"44",x"44",x"64",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"FF",x"FB",x"F5",x"F6",x"FF",x"FA",x"D1",x"FA",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"44",x"20",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"DB",x"FF",x"FF",x"FF",x"FF",x"F2",x"A4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"44",x"44",x"44",x"44",x"44",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"F5",x"FA",x"FF",x"FA",x"D1",x"FB",x"FF",x"F5",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"CC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"72",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"91",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"96",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"68",x"8C",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FB",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",
x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"92",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"64",x"AC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"F5",x"F6",x"F5",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"88",x"64",x"44",
x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"8C",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"88",x"64",x"44",x"44",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"BA",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"88",x"68",x"64",x"44",x"44",x"44",x"44",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F5",x"FA",x"FF",x"FF",x"FF",x"FB",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"CC",x"AC",x"88",x"68",x"64",x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"A4",x"F2",
x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"AC",x"AC",x"88",x"68",
x"68",x"64",x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C4",x"C4",
x"F6",x"FF",x"FF",x"FF",x"96",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"88",x"64",x"64",x"64",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"88",x"C4",x"C4",
x"C9",x"FB",x"FF",x"FF",x"96",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"CC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C4",x"C4",x"C4",
x"C4",x"E9",x"FF",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"88",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"96",x"C9",x"C4",x"C4",
x"C4",x"C4",x"F2",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D0",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D5",x"FF",x"FB",x"F5",x"FA",x"FF",x"FA",x"F5",x"FA",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FB",x"C5",x"C4",
x"C4",x"C4",x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"8C",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"FB",x"FA",x"D1",x"FA",x"FF",x"FA",x"D1",x"FA",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"F2",x"C4",
x"C4",x"C4",x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"96",x"FF",x"FF",x"FF",x"ED",
x"C4",x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"CC",x"AC",x"8C",x"64",x"44",x"64",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FF",x"FF",x"FF",x"FF",
x"C4",x"C4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"8C",x"88",
x"68",x"64",x"64",x"64",x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",
x"F6",x"68",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"F5",x"F5",x"FA",x"F5",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"8C",x"88",
x"68",x"64",x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"BA",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D0",x"AC",x"AC",x"AC",x"88",x"88",x"88",x"88",x"88",x"68",x"64",x"44",x"44",x"44",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"BA",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"44",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"BA",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FF",x"FF",x"FF",x"FF",x"FF",x"BA",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FF",x"FF",x"FF",x"FF",x"FF",x"96",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"FF",x"FF",x"FF",x"FF",x"DF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"88",x"88",x"88",x"88",x"88",
x"88",x"88",x"88",x"88",x"8C",x"8C",x"AC",x"AC",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FF",x"96",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"68",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"92",x"92",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D0",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"8C",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"44",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D0",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D0",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D0",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"44",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"8C",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",
x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",
x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"8C",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"64",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",
x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"64",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"64",x"CC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"64",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"64",x"44",x"44",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",
x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",x"CC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"64",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"68",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"68",x"AC",x"D1",x"D1",x"D1",
x"D1",x"AC",x"64",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",
x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"64",x"68",x"68",x"68",
x"64",x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",
x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",
x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",x"44",
x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",
x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"44",x"44",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"8C",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"88",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"68",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",x"44",
x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",x"44",
x"44",x"44",x"88",x"8C",x"8C",x"8C",x"88",x"68",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"44",x"44",x"44",x"44",x"40",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"24",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0");
	
	--Embbeded signals
	--Moving an object in the x axis
  signal x_axis  : integer range 0 to 640;
  
  --Offsets of all objects in screen
  signal offsetXC  : STD_LOGIC_VECTOR (9 downto 0);
  signal offsetYC  : STD_LOGIC_VECTOR (9 downto 0);
  
  --Addresses 
  signal Address : STD_LOGIC_VECTOR (16 downto 0);
  
  -- Definition of state names 
  type state_values is (front, left, right);
  signal pres_state, next_state: state_values;

  -- Data_In will be used to group input signals: Left, Right and Hazard
  signal   Data_In : std_logic_vector(1 downto 0);
  
begin

	-- Process which describes the "Current State Register"
  statereg: process (Clk, enable60, Rst)
  begin
    if (Rst='1') then 
      pres_state <= front;
    elsif (rising_edge(Clk) and enable60 = '1') then
      pres_state <= next_state;
    end if;
  end process statereg;
  
  -- Process that describes the "Next State Logic" section
  -- Group input signals for easier handling
  Data_In <= leftB & rightB;
  animation: process (pres_state, Data_In)
  begin
    case pres_state is
      when front => 
        case Data_In is
          when "10"   => next_state <= left;
          when "01"   => next_state <= right;
          when "00"   => next_state <= front;
          when others  => next_state <= front;
        end case;
        
      when right  => 
			case Data_In is
				 when "10"   => next_state <= front;
				 when "01"   => next_state <= right;
				 when "00"   => next_state <= front;
				 when others  => next_state <= front;
			  end case;
		
      when left => 
			case Data_In is
				 when "10"   => next_state <= left;
				 when "01"   => next_state <= front;
				 when "00"   => next_state <= front;
				 when others => next_state <= front;
			  end case;
      when others      => next_state <= front;
    end case;
  end process animation;
    
	--Calculates the address that will be taken from the memory for each object
  Address <= (Xin-offsetXC) + ((Yin-offsetYC)&"0000000");
  AddressCookie <= Address(13 downto 0);
  Address <= (Xin-offsetXC) + ((Yin-offsetYC)&"0000000");
  AddressCookieL <= Address(13 downto 0);
  Address <= (Xin-offsetXC) + ((Yin-offsetYC)&"0000000");
  AddressCookieR <= Address(13 downto 0);
  
  -- Process which describe the "Output Logic" section
  outputs: process (pres_state,AddressCookie,Color_Cookie)
  begin
    case pres_state is
      
      when front => Color_Cookie <= cookieF (conv_integer(AddressCookie ));
		when right => Color_Cookie <= cookieR (conv_integer(AddressCookieR));
		when left  => Color_Cookie <= cookieL (conv_integer(AddressCookieL));
      when others => null;
    end case;
  end process outputs;

 --The next process updates the cookie's positions according to the inputs from buttons
  Cookie: process (rightB, leftB, enable60,rst, x_axis, clk)
  begin
	 if (rst = '1') then
		 --Initial values (places cookie in the middle)
		 x_axis <= 256;
		 offsetYC <= CONV_STD_LOGIC_VECTOR(358, 10);
		 offsetXC <= CONV_STD_LOGIC_VECTOR(512, 10);
		 
	 elsif(rising_edge(clk)) then
		if(enable60 = '1') then
		 -- Updates the offset in X 
			offsetXC <= CONV_STD_LOGIC_VECTOR(640 - x_axis, 10);
			if (rightB = '1' and x_axis > 0) then
			-- Move to the right
				x_axis <= x_axis - 1;
			elsif (leftB = '1' and x_axis < 512) then
			-- Move to the left
				x_axis <= x_axis + 1;
			end if;
		end if;
	 end if;
  end process Cookie;
 
  -- Red Green Blue White
  process (En,Xin, Yin, AddressCookie, x_axis,Color_Cookie) 
  begin
    -- Check if pixel is in the active zone
	 if (En = '1') then
			--For drawing the cookie, we must check if the Xin and Yin are in the place the cookie will be drawn
			  if ((Xin>= (512 - x_axis) and Xin < (640 - x_axis)) and Yin > 352) then
				 Color <= Color_Cookie;
			  else
				 --In any other case, draw everything RED
				 Color <= "11100000"; -- RED
			  end if;
	 else
			-- Not in active zone, pixels should be OFF
			Color <= "00000000"; 
	 end if;
  end process;
  
    -- Send individual color to their channel
  R <= Color(7 downto 5);
  G <= Color(4 downto 2);
  B <= Color(1 downto 0);

end Behavioral;





