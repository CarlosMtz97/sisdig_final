----------------------------------------------------------------------------------
-- Company:      
-- Engineer:       
-- Create Date:     
-- Design Name: 
-- Module Name:    VGA_DISPLAY - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description:    
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
-- Commonly used libraries
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity VGA_DISPLAY is
  Generic
  ( n         : integer := 14;                    -- Number of Address bus lines, for an image of 128x128 pixels
	 m         : integer := 8);                    -- Number of Data bus lines
  port (
	 Xin       : in  STD_LOGIC_VECTOR(9 downto 0); -- Column screen coordinate
	 Yin       : in  STD_LOGIC_VECTOR(9 downto 0); -- Row screen coordinate
	 En        : in  STD_LOGIC;                    -- When '1', pixels can be drawn 
	 Enable60  : in  STD_LOGIC;                    -- Enable for cookie
	 rightB    : in  STD_LOGIC;                    -- Right button
	 leftB     : in  STD_LOGIC;                    -- Left button
	 rst       : in  STD_LOGIC;                    -- Reset
	 clk       : in  STD_LOGIC;                    -- Clock from FPGA
	 R   		  : out STD_LOGIC_VECTOR(2 downto 0); -- 3-bit Red channel
	 G   		  : out STD_LOGIC_VECTOR(2 downto 0); -- 3-bit Green channel
	 B   		  : out STD_LOGIC_VECTOR(1 downto 0));-- 2-bit Blue channel
end VGA_DISPLAY;


architecture Behavioral of VGA_DISPLAY is
  -- Embedded signal to group the colors into 1-byte
  -- The colors will be as follows:
  --  R2 R1 R0 G2 G1 G0 B1 B0
  signal Color : STD_LOGIC_VECTOR(7 downto 0); 
  
  --Addresses for the different images that will be displayed
  signal AddressCookie : STD_LOGIC_VECTOR(n-1 downto 0); --Super Cookie
  signal Data        : STD_LOGIC_VECTOR(m-1 downto 0);
  
  --Types of roms that will be used
  type objectImage is array (0 to (64**2) - 1) of STD_LOGIC_VECTOR (7 downto 0);
  type characterImage is array (0 to (128**2) - 1) of STD_LOGIC_VECTOR (7 downto 0);
  type kokoroImage is array (0 to (2**8) - 1) of STD_LOGIC_VECTOR (7 downto 0); --n=8 (8 bits) porque 2^n=2^8=256
 
  
  constant cookieS : characterImage := (
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FB",x"B2",x"8D",
x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"89",x"B1",x"DB",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"D6",x"8D",x"64",x"44",x"44",
x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"68",x"B2",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"DA",x"68",x"44",x"44",x"44",x"64",x"68",
x"88",x"8C",x"AC",x"AC",x"AD",x"AC",x"AC",x"AC",x"88",x"68",x"64",x"44",x"44",x"44",x"68",x"B2",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"8D",x"64",x"44",x"64",x"68",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"88",x"64",x"44",x"44",
x"68",x"DA",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",x"68",x"44",x"64",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"64",
x"44",x"64",x"B1",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"64",x"44",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"88",x"64",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"B2",x"64",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"64",x"44",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"B2",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"64",x"44",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"B6",x"64",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"89",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"DA",x"64",x"64",x"B1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",
x"F6",x"D1",x"D1",x"D1",x"D1",x"64",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"68",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",
x"FB",x"D1",x"D1",x"D1",x"D1",x"B1",x"64",x"44",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",
x"8D",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",
x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"64",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",
x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D5",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",
x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"F5",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FA",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",
x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"F5",x"FF",x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"D5",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"68",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",
x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"FF",x"FF",x"FA",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"64",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",
x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"68",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"68",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",
x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"D5",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"DB",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"AC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"8D",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"64",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"68",x"FF",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"68",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FF",x"FA",x"D5",x"FF",
x"FF",x"FB",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F5",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"DA",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FA",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"FF",
x"FF",x"FA",x"D5",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"F6",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B1",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"91",x"44",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D5",x"FA",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"FA",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"44",x"89",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"64",x"D1",x"D1",x"D1",
x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",
x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"68",x"D1",x"D1",x"D5",
x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"FA",x"FF",x"FF",x"FA",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",
x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"DB",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"44",x"88",x"D1",x"FB",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FA",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",
x"FF",x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"D6",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"8C",x"D1",x"FB",x"FF",
x"FB",x"FA",x"D5",x"D1",x"D1",x"D1",x"D5",x"F6",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"DF",
x"BB",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B2",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FA",x"D5",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"FF",x"F5",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"BB",x"13",
x"13",x"57",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B1",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D5",x"D1",
x"D1",x"D1",x"FF",x"F6",x"FF",x"D1",x"D1",x"FB",x"FA",x"D1",x"FF",x"FF",x"FF",x"9B",x"13",x"13",
x"13",x"13",x"9B",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AD",x"44",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FA",x"FA",x"FF",x"FA",x"FF",x"F5",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"77",x"13",x"13",x"13",
x"13",x"13",x"37",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FB",x"FF",x"9B",x"57",x"9B",x"DF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"F6",x"FF",x"F6",x"D1",x"F6",x"FF",x"FF",x"FF",x"57",x"13",x"13",x"13",x"13",
x"13",x"13",x"13",x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"DF",x"13",x"13",x"13",x"13",x"13",x"33",
x"77",x"FF",x"FF",x"D1",x"F6",x"D5",x"D1",x"D1",x"FA",x"FB",x"FF",x"33",x"13",x"13",x"13",x"13",
x"13",x"13",x"13",x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"77",x"13",x"13",x"13",x"13",x"13",x"13",
x"13",x"BF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"57",x"13",x"13",x"13",x"13",
x"13",x"13",x"57",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"91",x"44",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"37",x"13",x"13",x"13",x"13",x"13",x"13",
x"13",x"9B",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"BB",x"13",x"13",x"13",x"13",
x"13",x"13",x"DF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"57",x"13",x"13",x"13",x"13",x"13",x"13",
x"13",x"BB",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"77",x"13",x"13",x"13",
x"13",x"BB",x"FF",x"FF",x"F5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B1",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"9B",x"13",x"13",x"13",x"13",x"13",x"13",
x"13",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"DF",x"9B",x"9B",
x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B6",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",x"44",x"68",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C8",x"CC",x"D1",x"D1",x"FF",x"FF",x"33",x"13",x"13",x"13",x"13",x"13",
x"77",x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",
x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"D6",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"64",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C0",x"C4",x"D1",x"D1",x"FA",x"FF",x"DF",x"33",x"13",x"13",x"13",x"77",
x"FF",x"FF",x"D5",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"FB",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"44",x"AC",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C0",x"C0",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"BB",x"9B",x"DF",x"FF",
x"FF",x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"68",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"88",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C0",x"C0",x"CC",x"D1",x"D1",x"D1",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FA",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"8D",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"68",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"C4",x"C0",x"C4",x"D1",x"D1",x"D1",x"D1",x"D5",x"FA",x"FA",x"FA",x"D5",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"B2",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"64",x"B1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"CD",x"C0",x"C0",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"FB",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"88",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",x"C0",x"C0",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"68",x"FF",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"64",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"C8",x"C0",x"C0",x"C4",x"C8",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"B2",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"44",x"AC",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C4",x"C0",x"C0",x"C0",x"C4",x"C8",x"CC",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CD",x"CC",x"CD",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"68",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C4",x"C0",x"C0",x"C0",x"C0",x"C0",
x"C0",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C0",x"C0",x"C0",x"C0",x"C8",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"8D",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"44",
x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"CC",x"C8",x"C4",x"C4",
x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C4",x"C8",x"C8",x"CD",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",
x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"CD",x"CD",x"CD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",
x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",
x"64",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"B1",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"68",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"89",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"DA",x"B1",x"8D",x"8D",x"B2",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FF",x"68",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"68",x"64",x"44",x"44",x"44",x"44",x"64",x"B1",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"DB",x"64",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"88",x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"B1",x"64",x"44",x"68",x"B2",x"D6",x"D6",x"B1",x"64",x"44",x"8D",x"FF",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"DB",x"64",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"B1",x"44",x"64",x"D6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"89",x"44",x"8D",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"DB",x"68",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"64",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"D6",x"44",x"64",x"C0",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"68",x"44",
x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"B2",x"64",x"64",x"44",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",
x"64",x"64",x"64",x"8D",x"DB",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FF",x"68",x"64",x"C0",x"C0",x"C9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"64",
x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FB",x"89",x"44",x"64",x"AC",x"88",x"64",x"44",x"64",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",
x"88",x"D1",x"D1",x"88",x"64",x"B1",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"B2",x"44",x"A4",x"C0",x"C0",x"C0",x"ED",x"FB",x"D6",x"FF",x"FF",x"FB",x"F6",x"ED",x"84",
x"44",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"D6",x"64",x"44",x"68",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"AD",
x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"68",x"B6",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"68",x"68",x"C4",x"C0",x"C0",x"C0",x"84",x"64",x"44",x"64",x"A9",x"C0",x"C0",x"C0",x"C0",
x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",
x"8D",x"64",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"8D",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"DA",x"44",x"B2",x"F6",x"C0",x"C0",x"84",x"44",x"68",x"8D",x"64",x"64",x"C0",x"C0",x"C0",x"C0",
x"84",x"44",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"89",
x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"64",x"64",x"B2",x"FF",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"B1",x"64",x"DB",x"FF",x"F2",x"A0",x"64",x"68",x"FF",x"FF",x"D6",x"44",x"84",x"C0",x"C0",x"C0",
x"A0",x"64",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"68",x"44",
x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"8D",x"68",x"FF",x"FF",x"FF",x"B1",x"44",x"D6",x"E0",x"E0",x"FF",x"8D",x"64",x"C9",x"F6",x"FB",
x"FB",x"68",x"68",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"64",x"44",x"64",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FA",x"FA",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"64",x"D6",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"68",x"89",x"FF",x"FF",x"FF",x"8D",x"64",x"FF",x"E0",x"E0",x"E0",x"D6",x"44",x"B2",x"FF",x"FF",
x"FF",x"8D",x"64",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"B6",x"64",x"44",x"68",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",
x"D1",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"64",x"64",x"B2",x"FF",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"64",x"8D",x"FF",x"FF",x"FF",x"8D",x"68",x"FF",x"E0",x"E0",x"E0",x"FF",x"64",x"68",x"FF",x"FF",
x"FF",x"D6",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"B2",x"64",x"44",x"68",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"B1",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"64",x"8D",x"FF",x"FF",x"FF",x"8D",x"64",x"FF",x"E0",x"E0",x"FF",x"FF",x"8D",x"64",x"FF",x"FF",
x"FF",x"FB",x"64",x"B1",x"E0",x"E0",x"E0",x"E0",x"FF",x"B1",x"44",x"44",x"88",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",
x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"68",x"89",x"FF",x"FF",x"FF",x"D6",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"D6",x"FF",
x"FF",x"FF",x"68",x"68",x"E0",x"E0",x"E0",x"FF",x"8D",x"44",x"64",x"8C",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FB",x"FF",x"FA",x"FA",x"FF",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"B1",x"64",
x"64",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"8D",x"68",x"FF",x"FF",x"FF",x"FB",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"8D",x"FF",
x"FF",x"FF",x"8D",x"64",x"FF",x"E0",x"FF",x"8D",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"D1",x"FF",x"F5",x"F6",x"FF",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",
x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"B2",x"44",x"A4",x"C9",x"C4",x"C4",x"64",x"64",x"FF",x"E0",x"E0",x"E0",x"FF",x"68",x"68",x"FF",
x"FF",x"FF",x"B6",x"44",x"DA",x"FF",x"89",x"44",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FA",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"68",x"64",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"DB",x"64",x"84",x"C0",x"C0",x"C0",x"84",x"44",x"FB",x"E0",x"E0",x"E0",x"E0",x"91",x"64",x"FF",
x"FF",x"FF",x"FB",x"44",x"8D",x"68",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"FF",x"FF",x"FF",x"FB",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"64",x"D1",x"D1",x"AC",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"8C",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FF",x"68",x"64",x"A0",x"C0",x"C0",x"84",x"44",x"FF",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"A4",
x"C4",x"C9",x"F2",x"64",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FB",x"FB",x"FA",x"F6",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"AC",x"AC",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"DA",x"64",x"64",x"A4",x"84",x"64",x"68",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"84",
x"C0",x"C0",x"C0",x"64",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"64",x"88",x"64",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FF",x"B1",x"64",x"44",x"44",x"64",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"64",
x"C0",x"C0",x"C0",x"84",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"68",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"D6",x"91",x"B2",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"64",
x"C4",x"C0",x"C0",x"A0",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"68",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"D5",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"88",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"44",
x"D6",x"FF",x"FB",x"F2",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"8C",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",x"44",
x"B2",x"FF",x"FF",x"FF",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"8C",x"44",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"8D",x"44",
x"8D",x"FF",x"FF",x"FF",x"B1",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"44",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"68",x"44",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"64",x"44",
x"68",x"FF",x"FF",x"FF",x"D6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"B1",x"64",x"44",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"64",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"64",
x"64",x"FF",x"FF",x"FF",x"FB",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"F5",x"FF",x"D1",x"FA",x"FF",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",
x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"64",x"68",x"AC",
x"44",x"D6",x"FF",x"FF",x"FF",x"68",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"44",x"44",x"68",x"68",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FA",x"FA",x"F5",x"FF",x"FA",x"FF",x"FA",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",
x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",
x"44",x"B1",x"FF",x"FF",x"FF",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"68",x"44",x"64",x"B1",x"FF",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"FF",x"FF",x"FF",x"FF",x"FF",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",
x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"64",x"D1",x"D1",
x"64",x"89",x"FF",x"FF",x"FF",x"B2",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",
x"64",x"44",x"68",x"D6",x"E0",x"FB",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D5",x"FF",x"FF",x"FF",x"F6",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"44",
x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"88",x"D1",x"D1",
x"88",x"64",x"FF",x"FF",x"FF",x"DB",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"68",x"44",
x"44",x"8D",x"FF",x"E0",x"E0",x"D6",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"F5",x"F6",x"D5",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"68",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"AC",x"D1",x"D1",
x"8C",x"44",x"C9",x"E9",x"F2",x"F6",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"44",x"64",
x"B6",x"FF",x"E0",x"E0",x"E0",x"B2",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"64",x"DB",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"AC",x"D1",x"D1",
x"AC",x"44",x"A4",x"C0",x"C0",x"C0",x"64",x"64",x"D1",x"D1",x"AC",x"64",x"44",x"44",x"8D",x"FB",
x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"68",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"64",x"B6",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"AC",x"D1",x"D1",
x"D1",x"64",x"84",x"C0",x"C0",x"C0",x"84",x"44",x"AC",x"68",x"64",x"44",x"68",x"D6",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"68",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"AC",x"AC",x"8C",x"64",x"44",x"44",x"B2",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",x"44",x"68",x"D1",x"D1",
x"D1",x"68",x"64",x"C0",x"C0",x"C0",x"A4",x"44",x"44",x"44",x"64",x"B1",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"44",x"44",x"44",x"44",x"64",x"B6",x"FF",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"44",x"68",x"AC",
x"D1",x"88",x"64",x"CD",x"C9",x"C4",x"C0",x"64",x"64",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"FB",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"44",x"64",x"64",x"64",x"8D",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"64",x"44",x"44",
x"44",x"44",x"44",x"D6",x"FF",x"FF",x"F6",x"68",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"DA",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",x"D6",x"FB",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"8D",x"64",
x"64",x"64",x"44",x"B2",x"FF",x"FF",x"FF",x"8D",x"64",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"B6",x"44",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",
x"FB",x"DB",x"64",x"8D",x"FF",x"FF",x"FF",x"B6",x"44",x"DA",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"91",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"8D",x"64",x"FF",x"FF",x"FF",x"DB",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B2",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"B1",x"44",x"FB",x"FF",x"FF",x"FF",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"68",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"B1",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"D6",x"44",x"B6",x"FF",x"FF",x"FF",x"8D",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"64",x"8D",x"FF",x"FF",x"FF",x"B2",x"44",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FB",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"68",x"68",x"FF",x"FF",x"FF",x"DA",x"44",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"DA",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"8D",x"64",x"FF",x"FF",x"FF",x"FF",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"B6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"88",x"68",x"68",x"88",x"8C",x"AD",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"B6",x"44",x"D6",x"FF",x"FF",x"FF",x"68",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"B1",x"44",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"44",x"44",x"44",x"44",x"44",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FB",x"44",x"89",x"F2",x"FB",x"FF",x"B1",x"64",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"64",x"B6",x"D6",x"D6",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"64",x"64",x"C0",x"C0",x"C9",x"AD",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"88",x"68",x"FF",x"E0",x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"8D",x"64",x"C0",x"C0",x"C0",x"C0",x"64",x"B1",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"68",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"64",x"B1",x"E0",x"E0",x"E0",x"8D",x"44",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"89",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"A0",x"C0",x"C0",x"C0",x"64",x"68",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"44",x"DB",x"E0",x"E0",x"E0",x"8D",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"89",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"DA",x"44",x"A8",x"C9",x"C0",x"C0",x"84",x"64",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"DB",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"88",x"68",x"FF",x"E0",x"E0",x"E0",x"91",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"89",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"8D",x"FF",x"FF",x"F2",x"A4",x"44",x"DA",x"E0",x"E0",x"E0",
x"E0",x"E0",x"D6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"89",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"68",x"68",x"FF",x"FF",x"FF",x"DB",x"44",x"B2",x"E0",x"E0",x"E0",
x"E0",x"E0",x"B2",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"AC",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"89",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"B1",x"64",x"FB",x"FF",x"FF",x"FF",x"64",x"8D",x"E0",x"E0",x"E0",
x"E0",x"E0",x"8D",x"44",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"88",x"64",x"FF",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"D6",x"FF",x"FF",x"FF",x"8D",x"68",x"FF",x"E0",x"E0",
x"E0",x"E0",x"8D",x"44",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"B1",x"FF",x"FF",x"FF",x"B1",x"44",x"FB",x"E0",x"E0",
x"E0",x"FF",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"AC",x"64",x"B6",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"44",x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"68",x"FF",x"FF",x"FF",x"D6",x"44",x"B6",x"E0",x"E0",
x"E0",x"FF",x"64",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"88",x"64",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"64",x"FF",x"FF",x"FF",x"FF",x"44",x"8D",x"E0",x"E0",
x"E0",x"FB",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"B2",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B2",x"44",x"DB",x"FF",x"FF",x"FF",x"68",x"68",x"FF",x"E0",
x"E0",x"D6",x"44",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",
x"44",x"B1",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FB",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DA",x"44",x"B6",x"FF",x"FF",x"FF",x"8D",x"64",x"FF",x"E0",
x"E0",x"B6",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",
x"44",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"88",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"88",x"64",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"8D",x"FB",x"FF",x"FF",x"B6",x"44",x"DB",x"E0",
x"E0",x"B1",x"44",x"AC",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",
x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"68",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"68",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"64",x"C0",x"C4",x"ED",x"CD",x"44",x"D6",x"E0",
x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",
x"8D",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"91",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"91",x"64",x"C0",x"C0",x"C0",x"A0",x"44",x"B6",x"E0",
x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",
x"D6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"8D",x"64",x"AC",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"D6",x"44",x"84",x"C0",x"C0",x"A0",x"44",x"B6",x"E0",
x"E0",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",
x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"44",x"88",x"D1",x"D1",x"D1",x"D1",
x"D1",x"D1",x"D1",x"AC",x"44",x"8D",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"64",x"A0",x"C0",x"84",x"44",x"DB",x"E0",
x"E0",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"8D",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"64",x"64",x"AC",x"D1",x"D1",x"D1",
x"D1",x"D1",x"AC",x"64",x"64",x"DB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B6",x"44",x"64",x"64",x"44",x"68",x"FF",x"E0",
x"E0",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"8C",x"44",x"B6",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"B1",x"44",x"64",x"AD",x"D1",x"D1",
x"D1",x"8C",x"64",x"44",x"B2",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"B2",x"64",x"44",x"68",x"FF",x"E0",x"E0",
x"E0",x"68",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"FF",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"68",x"44",x"64",x"68",x"88",
x"64",x"44",x"44",x"B1",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",
x"E0",x"8D",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"8D",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",x"8D",x"64",x"44",x"44",
x"44",x"64",x"B6",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"91",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"68",x"64",x"DB",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"DB",x"B2",x"B1",
x"D6",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"D6",x"44",x"8C",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"AC",x"44",x"8D",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FF",x"64",x"64",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"D1",x"64",x"64",x"FB",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"B1",x"44",x"68",x"D1",x"D1",x"D1",x"D1",x"AC",x"64",x"64",x"D6",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FF",x"68",x"44",x"64",x"88",x"88",x"68",x"64",x"64",x"B6",x"FF",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FB",x"68",x"44",x"44",x"44",x"44",x"68",x"DA",x"FF",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"FF",x"B6",x"8D",x"8D",x"D6",x"FF",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0");
  

	--Embbeded signals
	--For moving an object in the x axis
  signal x_axis  : integer range 0 to 640;

  --Offsets of all objects in screen
  signal offsetXC  : STD_LOGIC_VECTOR (9 downto 0);
  signal offsetYC 
  : STD_LOGIC_VECTOR (9 downto 0);
  
  --Addresses that are used for making large operations
  signal Address : STD_LOGIC_VECTOR (16 downto 0);
  
begin

   --Calculates the address that will be taken from the memory for each object
  Address <= (Xin-offsetXC) + ((Yin-offsetYC)&"0000000");
  AddressCookie <= Address(13 downto 0);
  
 --The next process updates the cookie's positions according to the inputs from buttons
  Cookie: process (rightB, leftB, enable60,rst, x_axis, clk)
  begin
	 if (rst = '1') then
		--Initial values (places cookie in the middle)
		 x_axis <= 256;
		 offsetYC <= "0101100000";
		 offsetXC <= CONV_STD_LOGIC_VECTOR(512, 10);
	 elsif(rising_edge(clk)) then
		if(enable60 = '1') then
		 -- Updates the offset in Y 
			offsetXC <= CONV_STD_LOGIC_VECTOR(640 - x_axis, 10);
			if (rightB = '1' and x_axis > 0) then
			-- Move to the right
				x_axis <= x_axis - 1;
			elsif (leftB = '1' and x_axis < 512) then
			-- Move to the left
				x_axis <= x_axis + 1;
			end if;
		end if;
	 end if;
  end process Cookie;
  

  process (En,Xin, Yin, AddressCookie, x_axis) 
  begin
    -- Check if pixel is in the active zone
	 if (En = '1') then
			
			--For drawing the cookie, we must check if the Xin and Yin are in the place the cookie will be drawn
			  if ((Xin>= (512 - x_axis) and Xin < (640 - x_axis)) and Yin > 352) then
				 Color <= cookieS (conv_integer(AddressCookie));
			  else
				 --In any other case, draw everything RED
				 Color <= "11100000"; -- RED
			  end if;
	 else
			-- Not in active zone, pixels should be OFF
			Color <= "00000000"; 
	 end if;
  end process;
  
    -- Send individual color to their channel
  R <= Color(7 downto 5);
  G <= Color(4 downto 2);
  B <= Color(1 downto 0);

end Behavioral;





